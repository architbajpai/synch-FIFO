
class packet_fifo;
rand bit we,re;
rand bit [15:0] din;
bit [15:0] dout;
bit flagf,flage;

/*function void pre_randomize();
$display("we_pre:%0b	re_pre:%0b",we,re);
endfunction

function void post_randomize();
$display("we_post:%0b	re_post:%0b",we,re);
endfunction*/

/*task print();
$display("we=%b re=%b",we,re);
endtask*/

endclass


