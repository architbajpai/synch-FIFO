interface intf_fifo (input clk,rst);
bit we,re;
bit [15:0] din,dout;
bit flagf,flage;
endinterface